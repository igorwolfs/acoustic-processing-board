module top(
	