* Created by Paul Goedeke; July 10, 2018
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2018 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt TSV912 IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)

I_OS        ESDn MID 950F
I_B         25 MID 1P
V_GRp       60 MID 60
V_GRn       61 MID -60
V_ISCp      54 MID 54
V_ISCn      55 MID -54
V_ORn       34 VCLP -1.5
V11         59 33 0
V_ORp       32 VCLP 1.5
V12         58 31 0
V4          47 OUT 0
VCM_MIN     82 VEE_B -100M
VCM_MAX     83 VCC_B 100M
I_Q         VCC VEE 600U
V_OS        26 37 282.259U
C30         21 MID  3.18000000000000E-0016 
R69         MID 21   1MEG NOISELESS
G7          21 MID 22 MID  -1U
C29         22 MID 1.56F 
R80         MID 22   1MEG NOISELESS
G19         22 MID 23 MID  -1U
R51         ESDp 24   1M 
XVOS_VCM    25 26 VCC VEE VOS_SRC_0
S5          VEE ESDp VEE ESDp  S_VSWITCH_1
S4          VEE ESDn VEE ESDn  S_VSWITCH_2
S2          ESDn VCC ESDn VCC  S_VSWITCH_3
S3          ESDp VCC ESDp VCC  S_VSWITCH_4
C28         27 MID 1P 
R72         28 27   100 NOISELESS
C27         29 MID 1P 
R71         30 29   100 NOISELESS
R75         MID 31   1 NOISELESS
G14         31 MID 32 MID  -1
R74         33 MID   1 NOISELESS
G13         33 MID 34 MID  -1
R89         35 MID   1 NOISELESS
XVCCS_LIM_ZO 36 MID MID 35 VCCS_LIM_ZO_0
Xi_nn       ESDn MID FEMT_0
Xi_np       MID 37 FEMT_0
Xe_n        24 37 VNSE_0
C26         23 MID 3.18F 
R79         MID 23   1MEG NOISELESS
G18         23 MID VSENSE MID  -1U
C36         CLAMP MID 39.2N 
R68         MID CLAMP   1MEG NOISELESS
XVCCS_LIM_2 38 MID MID CLAMP VCCS_LIM_2_0
R44         MID 38   1MEG NOISELESS
XVCCS_LIM_1 39 40 MID 38 VCCS_LIM_1_0
R72_2       36 MID   1.11K NOISELESS
C31         36 41 15.92F 
R87         36 41   10K NOISELESS
R86         41 MID   1 NOISELESS
Gb1         41 MID 42 MID  -1
C22         43 MID 45F 
R85         42 43   10K NOISELESS
R84         42 44   90K NOISELESS
R83         44 MID   1 NOISELESS
G21         44 MID 45 MID  -6.5
C21         46 45 1.59U 
R55         45 MID   1.82K NOISELESS
R54         45 46   10K NOISELESS
Rdummy      MID 47   4K NOISELESS
Rx          47 35   40K NOISELESS
Rdc2        46 MID   1 NOISELESS
G10         46 MID CL_CLAMP 47  -60.61
R46         MID 48   3.572K NOISELESS
C14         48 49 15.9P 
R48         49 48   100MEG NOISELESS
G6          49 MID VEE_B MID  -99.34M
Rsrc1       MID 49   1 NOISELESS
R49         MID 50   3.572K NOISELESS
C16         50 51 15.9P 
R50         51 50   100MEG 
G9          51 MID VCC_B MID  -99.34M
Rsrc2       MID 51   1 NOISELESS
R81         MID 52   10.001K NOISELESS
C20         52 53 1.591P 
R82         53 52   100MEG NOISELESS
G20         53 MID ESDp MID  -100M
Rsrc3       MID 53   1 NOISELESS
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 2P 
XCL_AMP     54 55 VIMON MID 56 57 CLAMP_AMP_LO_0
S8          CLAMP 58 CLAMP 58  S_VSWITCH_5
S9          59 CLAMP 59 CLAMP  S_VSWITCH_6
XGR_AMP     60 61 62 MID 63 64 CLAMP_AMP_HI_0
R39         60 MID   1T NOISELESS
R37         61 MID   1T NOISELESS
R42         VSENSE 62   1M NOISELESS
C19         62 MID 1F 
R38         63 MID   1 NOISELESS
R36         MID 64   1 NOISELESS
R40         63 65   1M NOISELESS
R41         64 66   1M NOISELESS
C17         65 MID 1F 
C18         MID 66 1F 
XGR_SRC     65 66 CLAMP MID VCCS_LIM_GR_0
R21         56 MID   1 NOISELESS
R20         MID 57   1 NOISELESS
R29         56 67   1M NOISELESS
R30         57 68   1M NOISELESS
C9          67 MID 1F 
C8          MID 68 1F 
XCL_SRC     67 68 CL_CLAMP MID VCCS_LIM_4_0
R22         54 MID   1T NOISELESS
R19         MID 55   1T NOISELESS
XCLAWp      VIMON MID 69 VCC_B VCCS_LIM_CLAWP_0
XCLAWn      MID VIMON VEE_B 70 VCCS_LIM_CLAWN_0
R12         69 VCC_B   1K NOISELESS
R16         69 71   1M NOISELESS
R13         VEE_B 70   1K NOISELESS
R17         72 70   1M NOISELESS
C6          72 MID 1F 
C5          MID 71 1F 
G2          VCC_CLP MID 71 MID  -1M
R15         VCC_CLP MID   1K NOISELESS
G3          VEE_CLP MID 72 MID  -1M
R14         MID VEE_CLP   1K NOISELESS
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 73 74 CLAMP_AMP_LO_0
R26         VCC_CLP MID   1T NOISELESS
R23         VEE_CLP MID   1T NOISELESS
R25         73 MID   1 NOISELESS
R24         MID 74   1 NOISELESS
R27         73 75   1M NOISELESS
R28         74 76   1M NOISELESS
C11         75 MID 1F 
C10         MID 76 1F 
XCLAW_SRC   75 76 CLAW_CLAMP MID VCCS_LIM_3_0
H2          30 MID V11 -1
H3          28 MID V12 1
C12         SW_OL MID 1N 
R32         77 SW_OL   100 NOISELESS
R31         77 MID   1 NOISELESS
XOL_SENSE   MID 77 29 27 OL_SENSE_0
S1          46 45 SW_OL MID  S_VSWITCH_7
H1          78 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_8
S6          OUT VCC OUT VCC  S_VSWITCH_9
R11         MID 79   1T NOISELESS
R18         79 VOUT_S   100 NOISELESS
C7          VOUT_S MID 1P 
E5          79 MID OUT MID  1
C13         VIMON MID 10P 
R33         78 VIMON   100 NOISELESS
R10         MID 78   1T NOISELESS
R47         80 VCLP   100 NOISELESS
C24         VCLP MID 100P 
E4          80 MID CL_CLAMP MID  1
R62         MID CL_CLAMP   1K NOISELESS
G4          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP   1K NOISELESS
G8          CLAW_CLAMP MID 21 MID  -1M
R43         MID VSENSE   1K NOISELESS
G15         VSENSE MID CLAMP MID  -1M
C4          39 MID 1F 
R9          39 81   1M NOISELESS
R7          MID 82   1T NOISELESS
R6          83 MID   1T NOISELESS
R8          MID 81   1 NOISELESS
XVCM_CLAMP  84 MID 81 MID 83 82 VCCS_EXT_LIM_0
E1          MID 0 85 0  1
R77         VEE_B 0   1 NOISELESS
R5          86 VEE_B   1M NOISELESS
C3          86 0 1F 
R60         85 86   1MEG NOISELESS
C1          85 0 1 
R3          85 0   1T NOISELESS
R59         87 85   1MEG NOISELESS
C2          87 0 1F 
R4          VCC_B 87   1M NOISELESS
R76         VCC_B 0   1 NOISELESS
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R67         88 84   1K NOISELESS
G1          84 88 50 48  -1M
R2          40 ESDn   1M NOISELESS
R1          88 89   1M NOISELESS
R58         25 89   1K NOISELESS
G5          89 25 52 MID  -1M
C_CMn       ESDn MID 4P 
C_CMp       MID ESDp 4P 
R53         ESDn MID   1T NOISELESS
R52         MID ESDp   1T NOISELESS
R35         IN- ESDn   10M NOISELESS
R34         IN+ ESDp   10M NOISELESS

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_8 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_9 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)

.ENDS TSV912
*
.SUBCKT VOS_SRC_0  V+ V- REF+ REF-
E1 V+ 1 TABLE {(V(REF+, V-))} =
+(0, 1.6E-3)
+(1, 1.6E-3)
+(1.3, 0)
+(5.5, 0)
E2 1 V- TABLE {(V(V-, REF-))}=
+(-0.7, -2E-4)
+(-0.5, -2E-4)
+(-0.4, 0)
+(5.5, 0)
.ENDS VOS_SRC_0 
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 10
.PARAM IPOS = 10E3
.PARAM INEG = -10E3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=7
.PARAM NVRF=7
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16 cjo=.1f
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS FEMT_0 
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=10
.PARAM NLF=100
.PARAM NVR=11
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16 cjo=.1f
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS VNSE_0 
*


.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 24.63E-3
.PARAM IPOS = 0.247
.PARAM INEG = -0.247
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.494
.PARAM INEG = -0.494
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.228
.PARAM INEG = -0.228
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAWP_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 5E-5)
+(10, 1.38E-4 )
+(20, 2.93E-4)
+(30, 4.78E-4)
+(40, 7.21E-4)
+(45, 8.95E-4)
+(47, 9.92E-4)
+(50, 1.24E-3)
+(52, 1.59E-3)
+(54, 2.23E-3)
.ENDS VCCS_LIM_CLAWP_0 
*


.SUBCKT VCCS_LIM_CLAWN_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 5E-5 )
+(10, 1.29E-4)
+(20, 2.77E-4)
+(30, 4.52E-4)
+(40, 6.77E-4)
+(45, 8.31E-4)
+(47, 9.09E-4)
+(50, 1.08E-3)
+(52, 1.3E-3)
+(54, 2.25E-3)
.ENDS VCCS_LIM_CLAWN_0 
*


.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.114
.PARAM INEG = -0.114
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIM_3_0 
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*


