* OPA2991 - Rev. A
* Created by Bala Ravi; September 09, 2019
* Created with Green-Williams-Lis Op Amp Macro-model Architecture
* Copyright 2019 by Texas Instruments Corporation
******************************************************
* MACRO-MODEL SIMULATED PARAMETERS:
******************************************************
* OPEN-LOOP GAIN AND PHASE VS. FREQUENCY  WITH RL, CL EFFECTS (Aol)
* UNITY GAIN BANDWIDTH (GBW)
* INPUT COMMON-MODE REJECTION RATIO VS. FREQUENCY (CMRR)
* POWER SUPPLY REJECTION RATIO VS. FREQUENCY (PSRR)
* DIFFERENTIAL INPUT IMPEDANCE (Zid)
* COMMON-MODE INPUT IMPEDANCE (Zic)
* OPEN-LOOP OUTPUT IMPEDANCE VS. FREQUENCY (Zo)
* OUTPUT CURRENT THROUGH THE SUPPLY (Iout)
* INPUT VOLTAGE NOISE DENSITY VS. FREQUENCY (en)
* INPUT CURRENT NOISE DENSITY VS. FREQUENCY (in)
* OUTPUT VOLTAGE SWING vs. OUTPUT CURRENT (Vo)
* SHORT-CIRCUIT OUTPUT CURRENT (Isc)
* QUIESCENT CURRENT (Iq)
* SETTLING TIME VS. CAPACITIVE LOAD (ts)
* SLEW RATE (SR)
* SMALL SIGNAL OVERSHOOT VS. CAPACITIVE LOAD
* LARGE SIGNAL RESPONSE
* OVERLOAD RECOVERY TIME (tor)
* INPUT BIAS CURRENT (Ib)
* INPUT OFFSET CURRENT (Ios)
* INPUT OFFSET VOLTAGE (Vos)
* INPUT COMMON-MODE VOLTAGE RANGE (Vcm)
* INPUT OFFSET VOLTAGE VS. INPUT COMMON-MODE VOLTAGE (Vos vs. Vcm)
* INPUT/OUTPUT ESD CELLS (ESDin, ESDout)
******************************************************
.subckt OPA2991 IN+ IN- VCC VEE OUT
******************************************************
* MODEL DEFINITIONS:
.model BB_SW VSWITCH(Ron=50 Roff=1e12 Von=700e-3 Voff=0)
.model ESD_SW VSWITCH(Ron=50 Roff=1e12 Von=250e-3 Voff=0)
.model OL_SW VSWITCH(Ron=1e-3 Roff=1e9 Von=900e-3 Voff=800e-3)
.model OR_SW VSWITCH(Ron=10e-3 Roff=1e9 Von=1e-3 Voff=0)
.model R_NOISELESS RES(T_ABS=-273.15)
******************************************************

VS1         25 26 124.96U
I_OS        ESDn MID 0
I_B         26 MID 10P
V_GRp       56 MID 110
V_GRn       57 MID -110
V_ISCp      50 MID 80
V_ISCn      51 MID -80
V_ORn       34 VCLP -12
V11         55 33 0
V_ORp       32 VCLP 12
V12         54 31 0
V4          43 OUT 0
VCM_MIN     78 VEE_B -200M
VCM_MAX     79 VCC_B 200M
I_Q         VCC VEE 560U
GVCCS4      22 MID 21 MID  -1
R64         23 MID R_NOISELESS 1 
C22         24 MID 159F  
R63         21 24 R_NOISELESS 10K 
R62         23 21 R_NOISELESS 37.6K 
XIn11       ESDn MID FEMT_0
Xi_n        MID 26 FEMT_0
Xe_n        ESDp 26 VNSE_0
S5          VEE ESDp VEE ESDp  S_VSWITCH_1
S4          VEE ESDn VEE ESDn  S_VSWITCH_2
S2          ESDn VCC ESDn VCC  S_VSWITCH_3
S3          ESDp VCC ESDp VCC  S_VSWITCH_4
C28         27 MID 1P  
R77         28 27 R_NOISELESS 100 
C27         29 MID 1P  
R76         30 29 R_NOISELESS 100 
R75         MID 31 R_NOISELESS 1 
GVCCS8      31 MID 32 MID  -1
R74         33 MID R_NOISELESS 1 
GVCCS7      33 MID 34 MID  -1
R73         35 MID R_NOISELESS 1 
XVCCS_LIM_ZO 36 MID MID 35 VCCS_LIM_ZO_0
C25         37 MID 53.05F  
R69         MID 37 R_NOISELESS 1MEG 
GVCCS6      37 MID VSENSE MID  -1U
C20         CLAMP MID 289.4N  
R68         MID CLAMP R_NOISELESS 1MEG 
XVCCS_LIM_2 38 MID MID CLAMP VCCS_LIM_2_0
R44         MID 38 R_NOISELESS 1MEG 
XVCCS_LIM_1 39 40 MID 38 VCCS_LIM_1_0
R72         36 MID R_NOISELESS 2.5 
C26         36 22 636.6F  
R71         36 22 R_NOISELESS 10K 
R70         22 MID R_NOISELESS 1 
GVCCS3      23 MID 41 MID  -8.5
C21         42 41 22.3P  
R51         41 MID R_NOISELESS 3.51K 
R50         41 42 R_NOISELESS 10K 
Rdummy      MID 43 R_NOISELESS 7.97K 
Rx          43 35 R_NOISELESS 79.7K 
Rdc         42 MID R_NOISELESS 1 
G_Aol_Zo    42 MID CL_CLAMP 43  -40
R61         MID 44 R_NOISELESS 2 
C16         44 45 3.98N  
R58         45 44 R_NOISELESS 100MEG 
GVCCS2      45 MID VEE_B MID  -1.81
R57         MID 45 R_NOISELESS 1 
R56         MID 46 R_NOISELESS 2 
C15         46 47 3.98N  
R55         47 46 R_NOISELESS 100MEG 
GVCCS1      47 MID VCC_B MID  -1.81
R54         MID 47 R_NOISELESS 1 
R49         MID 48 R_NOISELESS 2K 
C14         48 49 198.9P  
R48         49 48 R_NOISELESS 100MEG 
G_adjust    49 MID ESDp MID  -60.53M
Rsrc        MID 49 R_NOISELESS 1 
XIQPos      VIMON MID MID VCC VCCS_LIMIT_IQ_0
XIQNeg      MID VIMON VEE MID VCCS_LIMIT_IQ_0
C_DIFF      ESDp ESDn 3P  
XCL_AMP     50 51 VIMON MID 52 53 CLAMP_AMP_LO_0
SOR_SWp     CLAMP 54 CLAMP 54  S_VSWITCH_5
SOR_SWn     55 CLAMP 55 CLAMP  S_VSWITCH_6
XGR_AMP     56 57 58 MID 59 60 CLAMP_AMP_HI_0
R39         56 MID R_NOISELESS 1T 
R37         57 MID R_NOISELESS 1T 
R42         VSENSE 58 R_NOISELESS 1M 
C19         58 MID 1F  
R38         59 MID R_NOISELESS 1 
R36         MID 60 R_NOISELESS 1 
R40         59 61 R_NOISELESS 1M 
R41         60 62 R_NOISELESS 1M 
C17         61 MID 1F  
C18         MID 62 1F  
XGR_SRC     61 62 CLAMP MID VCCS_LIM_GR_0
R21         52 MID R_NOISELESS 1 
R20         MID 53 R_NOISELESS 1 
R29         52 63 R_NOISELESS 1M 
R30         53 64 R_NOISELESS 1M 
C9          63 MID 1F  
C8          MID 64 1F  
XCL_SRC     63 64 CL_CLAMP MID VCCS_LIM_4_0
R22         50 MID R_NOISELESS 1T 
R19         MID 51 R_NOISELESS 1T 
XCLAWp      VIMON MID 65 VCC_B VCCS_LIM_CLAW+_0
XCLAWn      MID VIMON VEE_B 66 VCCS_LIM_CLAW-_0
R12         65 VCC_B R_NOISELESS 1K 
R16         65 67 R_NOISELESS 1M 
R13         VEE_B 66 R_NOISELESS 1K 
R17         68 66 R_NOISELESS 1M 
C6          68 MID 1F  
C5          MID 67 1F  
G2          VCC_CLP MID 67 MID  -1M
R15         VCC_CLP MID R_NOISELESS 1K 
G3          VEE_CLP MID 68 MID  -1M
R14         MID VEE_CLP R_NOISELESS 1K 
XCLAW_AMP   VCC_CLP VEE_CLP VOUT_S MID 69 70 CLAMP_AMP_LO_0
R26         VCC_CLP MID R_NOISELESS 1T 
R23         VEE_CLP MID R_NOISELESS 1T 
R25         69 MID R_NOISELESS 1 
R24         MID 70 R_NOISELESS 1 
R27         69 71 R_NOISELESS 1M 
R28         70 72 R_NOISELESS 1M 
C11         71 MID 1F  
C10         MID 72 1F  
XCLAW_SRC   71 72 CLAW_CLAMP MID VCCS_LIM_3_0
H2          30 MID V11 -1
H3          28 MID V12 1
C12         SW_OL MID 100P  
R32         73 SW_OL R_NOISELESS 100 
R31         73 MID R_NOISELESS 1 
XOL_SENSE   MID 73 29 27 OL_SENSE_0
S1          42 41 SW_OL MID  S_VSWITCH_7
H1          74 MID V4 1K
S7          VEE OUT VEE OUT  S_VSWITCH_8
S6          OUT VCC OUT VCC  S_VSWITCH_9
R11         MID 75 R_NOISELESS 1T 
R18         75 VOUT_S R_NOISELESS 100 
C7          VOUT_S MID 1N  
E5          75 MID OUT MID  1
C13         VIMON MID 1N  
R33         74 VIMON R_NOISELESS 100 
R10         MID 74 R_NOISELESS 1T 
R47         76 VCLP R_NOISELESS 100 
C24         VCLP MID 100P  
E4          76 MID CL_CLAMP MID  1
R46         MID CL_CLAMP R_NOISELESS 1K 
G9          CL_CLAMP MID CLAW_CLAMP MID  -1M
R45         MID CLAW_CLAMP R_NOISELESS 1K 
G8          CLAW_CLAMP MID 37 MID  -1M
R43         MID VSENSE R_NOISELESS 1K 
G15         VSENSE MID CLAMP MID  -1M
C4          39 MID 1F  
R9          39 77 R_NOISELESS 1M 
R7          MID 78 R_NOISELESS 1T 
R6          79 MID R_NOISELESS 1T 
R8          MID 77 R_NOISELESS 1 
XVCM_CLAMP  80 MID 77 MID 79 78 VCCS_EXT_LIM_0
E1          MID 0 81 0  1
R89         VEE_B 0 R_NOISELESS 1 
R5          82 VEE_B R_NOISELESS 1M 
C3          82 0 1F  
R60         81 82 R_NOISELESS 1MEG 
C1          81 0 1  
R3          81 0 R_NOISELESS 1T 
R59         83 81 R_NOISELESS 1MEG 
C2          83 0 1F  
R4          VCC_B 83 R_NOISELESS 1M 
R88         VCC_B 0 R_NOISELESS 1 
G17         VEE_B 0 VEE 0  -1
G16         VCC_B 0 VCC 0  -1
R_PSR       84 80 R_NOISELESS 1K 
G_PSR       80 84 46 44  -1M
R2          40 ESDn R_NOISELESS 1M 
R1          84 85 R_NOISELESS 1M 
R_CMR       25 85 R_NOISELESS 1K 
G_CMR       85 25 48 MID  -1M
C_CMn       ESDn MID 1P  
C_CMp       MID ESDp 1P  
R53         ESDn MID R_NOISELESS 1T 
R52         MID ESDp R_NOISELESS 1T 
R35         IN- ESDn R_NOISELESS 10M 
R34         IN+ ESDp R_NOISELESS 10M 

.MODEL S_VSWITCH_1 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=1T VON=10M VOFF=0)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_8 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)
.MODEL S_VSWITCH_9 VSWITCH (RON=50 ROFF=1T VON=500M VOFF=100M)

.ENDS OPA2991
*
.SUBCKT FEMT_0  1 2
.PARAM FLWF=1E-3
.PARAM NLFF=2
.PARAM NVRF=2
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
.ENDS
*


.SUBCKT VNSE_0  1 2
.PARAM FLW=0.1
.PARAM NLF=340
.PARAM NVR=9.39
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
.ENDS
*


.SUBCKT VCCS_LIM_ZO_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 4E3
.PARAM IPOS = 50E3
.PARAM INEG = -50E3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_2_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 8.577E-2
.PARAM IPOS = 5.788
.PARAM INEG = -5.788
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_1_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-4
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIMIT_IQ_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1E-3
G1 IOUT- IOUT+ VALUE={IF( (V(VC+,VC-)<=0),0,GAIN*V(VC+,VC-) )}
.ENDS
*


.SUBCKT CLAMP_AMP_LO_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=1
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT CLAMP_AMP_HI_0  VC+ VC- VIN COM VO+ VO-
.PARAM G=10
GVO+ COM VO+ VALUE = {IF(V(VIN,COM)>V(VC+,COM),((V(VIN,COM)-V(VC+,COM))*G),0)}
GVO- COM VO- VALUE = {IF(V(VIN,COM)<V(VC-,COM),((V(VC-,COM)-V(VIN,COM))*G),0)}
.ENDS
*


.SUBCKT VCCS_LIM_GR_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 0.0276
.PARAM INEG = -0.04416
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_4_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 12
.PARAM INEG = -12
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT VCCS_LIM_CLAW+_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1.00E-5)
+(30, 6.2E-4)
+(40, 8.6E-4)
+(60, 1.45E-3)
+(80, 2.5E-3)
+(83, 2.97E-3)
+(84.5, 4.03E-2)
.ENDS 
*


.SUBCKT VCCS_LIM_CLAW-_0  VC+ VC- IOUT+ IOUT-
G1 IOUT+ IOUT- TABLE {ABS(V(VC+,VC-))} =
+(0, 1E-5)
+(50, 9.8E-4)
+(60, 1.26E-3)
+(80, 2.19E-3)
+(82, 2.47E-3)
+(83, 2.72E-3)
+(84.45, 1.92E-2)
.ENDS
*



.SUBCKT VCCS_LIM_3_0  VC+ VC- IOUT+ IOUT-
.PARAM GAIN = 1
.PARAM IPOS = 550E-3
.PARAM INEG = -550E-3
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS
*


.SUBCKT OL_SENSE_0  COM SW+ OLN  OLP
GSW+ COM SW+ VALUE = {IF((V(OLN,COM)>10E-3 | V(OLP,COM)>10E-3),1,0)}
.ENDS
*


.SUBCKT VCCS_EXT_LIM_0  VIN+ VIN- IOUT- IOUT+ VP+ VP-
.PARAM GAIN = 1
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VIN+,VIN-),V(VP-,VIN-), V(VP+,VIN-))}
.ENDS
*


