module testbench;
	reg 