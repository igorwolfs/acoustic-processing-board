`timescale 1ns / 1ps

//
// RGMII Functional Interface Driver (Lattice ECP5 Verilog)
//
// This module provides a functional RGMII interface, converting the DDR PHY
// signals to a simpler, SDR application interface within the FPGA. This version
// is specifically adapted for Lattice ECP5 FPGAs.
//
// It uses IDDRX1F and ODDRX1F primitives to manage the double-data-rate conversion.
//
module rgmii (
    // --- System Inputs ---
    input        RESET_N,        // Active-low reset

    // --- Application Interface (SDR) ---
    output [7:0] RX_DATA,        // Received data byte
    output       RX_DV,          // Received data valid
    input  [7:0] TX_DATA,        // Transmit data byte
    input        TX_DV,          // Transmit data valid

    // --- RGMII PHY Interface (DDR) ---
    input        RGMII_RX_CLK,   // 125 MHz clock from PHY
    input        RGMII_RX_CTL,   // Contains RX_DV
    input  [3:0] RGMII_RX_D,

    output       RGMII_TX_CLK,   // 125 MHz clock to PHY
    output       RGMII_TX_CTL,   // Contains TX_EN
    output [3:0] RGMII_TX_D,

    // Management Interface (Stubbed)
    input        MDIO_CLK,
    inout        MDIO_DATA
);

    // --- Clocking ---
    // For Lattice ECP5, the synthesis tool infers the global clock buffer.
    // There is no need to instantiate a CLKBUF primitive. The tool will
    // automatically place RGMII_RX_CLK on a global clock network if it is
    // connected to a PCLK pin and/or drives many loads.
    //
    // It is critical to add a frequency constraint to your .lpf file, for example:
    // FREQUENCY PORT "RGMII_RX_CLK" 125.0 MHz;

    // In a real design, RGMII_TX_CLK should be generated by a PLL, phase-aligned
    // with RGMII_RX_CLK. For this example, we forward the RX clock.
    assign RGMII_TX_CLK = RGMII_RX_CLK;


    // --- RX Path (PHY -> FPGA Application) ---
    // Deserialize the DDR RGMII input to an 8-bit SDR bus for the application.
    wire rx_ctl_sdr;
    wire [7:0] rx_data_sdr;
    wire rst_sync = !RESET_N; // ECP5 primitives use active-high reset

    // Capture RX_CTL (Data Valid) signal using an IDDRX1F primitive.
    IDDRX1F iddrx1f_rx_ctl (
        .D(RGMII_RX_CTL),
        .SCLK(RGMII_RX_CLK), // Clocked directly by the input clock
        .RST(rst_sync),
        .Q0(rx_ctl_sdr), // Data from rising edge
        .Q1()           // Data from falling edge (unused for RX_CTL)
    );

    // Capture the 4-bit DDR data bus into an 8-bit SDR register.
    genvar i;
    generate
        for (i = 0; i < 4; i = i + 1) begin : gen_iddr_rx
            IDDRX1F iddrx1f_rx_data (
                .D(RGMII_RX_D[i]),
                .SCLK(RGMII_RX_CLK), // Clocked directly by the input clock
                .RST(rst_sync),
                .Q0(rx_data_sdr[i]),   // Rising edge data
                .Q1(rx_data_sdr[i+4])  // Falling edge data
            );
        end
    endgenerate

    // Assign deserialized signals to the application interface
    assign RX_DV   = rx_ctl_sdr;
    assign RX_DATA = rx_data_sdr;


    // --- TX Path (FPGA Application -> PHY) ---
    // Serialize the 8-bit SDR data from the application to the DDR RGMII output.
    
    // Drive TX_CTL (Transmit Enable) using an ODDRX1F primitive.
    ODDRX1F oddrx1f_tx_ctl (
        .D0(TX_DV),       // Data for rising edge
        .D1(TX_DV),       // Data for falling edge
        .SCLK(RGMII_TX_CLK),
        .RST(rst_sync),
        .Q(RGMII_TX_CTL)
    );

    // Drive the 4-bit DDR data bus from the 8-bit SDR application data.
    generate
        for (i = 0; i < 4; i = i + 1) begin : gen_oddr_tx
            ODDRX1F oddrx1f_tx_data (
                .D0(TX_DATA[i]),   // Lower nibble on rising edge
                .D1(TX_DATA[i+4]), // Upper nibble on falling edge
                .SCLK(RGMII_TX_CLK),
                .RST(rst_sync),
                .Q(RGMII_TX_D[i])
            );
        end
    endgenerate


    // --- MDIO Interface Stub ---
    // Assign to high-impedance as we are not implementing MDIO logic.
    assign MDIO_DATA = 1'bz;

endmodule