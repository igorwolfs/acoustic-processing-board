.SUBCKT irf740lc 1 2 3
* Model generated on Aug 17, 98
* MODEL FORMAT: SPICE3
* Symmetry POWER MOS Model (Version 1.0)
* External Node Designations
* Node 1 -> Drain
* Node 2 -> Gate
* Node 3 -> Source
M1 9 7 8 8 MM L=100u W=100u
.MODEL MM NMOS LEVEL=1 IS=1e-32
+VTO=4 LAMBDA=0 KP=1.5638
+CGSO=1.09984e-05 CGDO=1e-11
RS 8 3 0.0001
D1 3 1 MD
.MODEL MD D IS=2.35458e-11 RS=0.0192633 N=1.11352 BV=400
+IBV=0.00025 EG=1 XTI=3.06659 TT=0
+CJO=1.69617e-09 VJ=2.25185 M=0.9 FC=0.5
RDS 3 1 1e+06
RD 9 1 0.401573
RG 2 7 5.55712
D2 4 5 MD1
.MODEL MD1 D IS=1e-32 N=50
+CJO=1.15293e-09 VJ=0.840745 M=0.9 FC=1e-08
D3 0 5 MD2
.MODEL MD2 D IS=1e-10 N=0.573951 RS=3e-06
RL 5 10 1
FI2 7 9 VFI2 -1
VFI2 4 0 0
EV16 10 0 9 7 1
CAP 11 10 1.15293e-09
FI1 7 9 VFI1 -1
VFI1 11 6 0
RCAP 6 10 1
D4 0 6 MD3
.MODEL MD3 D IS=1e-10 N=0.573951
.ENDS irf740lc
